library verilog;
use verilog.vl_types.all;
entity TRCUTtb is
end TRCUTtb;
