`timescale 1ns/1ps

module LFSR16_18211(
  input clk,
  output reg [15:0] LFSR = 65535
);

wire feedback = LFSR[15];

always @(posedge clk)
begin
  LFSR[0] <= feedback;
  LFSR[1] <= LFSR[0];
  LFSR[2] <= LFSR[1];
  LFSR[3] <= LFSR[2];
  LFSR[4] <= LFSR[3] ^ feedback;
  LFSR[5] <= LFSR[4];
  LFSR[6] <= LFSR[5];
  LFSR[7] <= LFSR[6];
  LFSR[8] <= LFSR[7];
  LFSR[9] <= LFSR[8] ^ feedback;
  LFSR[10] <= LFSR[9];
  LFSR[11] <= LFSR[10];
  LFSR[12] <= LFSR[11];
  LFSR[13] <= LFSR[12];
  LFSR[14] <= LFSR[13];
  LFSR[15] <= LFSR[14] ^ feedback;
end
endmodule
