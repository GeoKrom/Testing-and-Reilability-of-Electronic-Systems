library verilog;
use verilog.vl_types.all;
entity TRCUTwithMISRtb is
end TRCUTwithMISRtb;
