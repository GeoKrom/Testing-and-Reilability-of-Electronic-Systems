library verilog;
use verilog.vl_types.all;
entity SDFFChaintb is
end SDFFChaintb;
